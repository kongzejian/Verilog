`timescale 1ns/1ns

module wire0(
    input in0,
    output out1
);
assign out1=in0;
endmodule
