`timescale 1ns/1ns

module top_module(
    input a,b,
    output x,y,z
);
assign z=a;
assign x=b;
assign y=b;
endmodule
