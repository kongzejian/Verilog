`timescale 1ns/1ns

module top_module( 
    input a, 
    input b, 
    output c );
    assign c=a^b;

endmodule
