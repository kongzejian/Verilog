`timescale 1ns/1ns
module top_module( 
    input a, 
    input b, 
    input c,
    output d );
assign d=a&b&c;
    
endmodule
